`timescale 1ns / 1ps

module tb_alu;

  logic [15:0] x;
  logic [15:0] y;
  bit   zx;    /* zero   x */
  bit   nx;    /* negate x */
  bit   zy;    /* zero   y */
  bit   ny;    /* negate y */
  bit   f;     /* 0: and, 1: add */
  bit   no;    /* negate output */
  logic [15:0] out;
  bit   zr;    /* output is zero */
  bit   ng;    /* output is negative */

  typedef struct packed {
    logic [15:0] x;
    logic [15:0] y;
    bit zx;
    bit nx;
    bit zy;
    bit ny;
    bit f;
    bit no;
  } tc_in_t;

  typedef struct packed {
    tc_in_t in;
    logic [15:0] out;
    bit zr;
    bit ng;
  } test_case_t;

  /* verilog_lint: waive-start line-length */
  /* verilog_format: off */
  test_case_t test_cases[] = '{
  /* x                    y                     zx    nx    zy    ny    f     no    out                   zr    ng   */
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 16'b0000000000000000, 1'b1, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 16'b0000000000000001, 1'b0, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 16'b0000000000000000, 1'b1, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 16'b0000000000000000, 1'b1, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 16'b0000000000000000, 1'b1, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 16'b0000000000000001, 1'b0, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 16'b0000000000000001, 1'b0, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 16'b0000000000000000, 1'b1, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 16'b1111111111111110, 1'b0, 1'b1 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 16'b0000000000000001, 1'b0, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 16'b0000000000000000, 1'b1, 1'b0 },
  { 16'b0000000000000000, 16'b1111111111111111, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 16'b0000000000000000, 1'b1, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 16'b0000000000000001, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 16'b1111111111111111, 1'b0, 1'b1 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 16'b0000000000010001, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 16'b0000000000000011, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 16'b1111111111101110, 1'b0, 1'b1 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 16'b1111111111111100, 1'b0, 1'b1 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 16'b1111111111101111, 1'b0, 1'b1 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 16'b1111111111111101, 1'b0, 1'b1 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 16'b0000000000010010, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 16'b0000000000000100, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 16'b0000000000010000, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 16'b0000000000000010, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 16'b0000000000010100, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 16'b0000000000001110, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 16'b1111111111110010, 1'b0, 1'b1 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 16'b0000000000000001, 1'b0, 1'b0 },
  { 16'b0000000000010001, 16'b0000000000000011, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 16'b0000000000010011, 1'b0, 1'b0 }
};
  /* verilog_lint: waive-end line-length */
  /* verilog_format: on */

  alu dut (.*);

  initial begin
    foreach (test_cases[i]) begin
      {x, y, zx, nx, zy, ny, f, no} = test_cases[i].in;
      #10;
      $monitor("@%0t: x=%h y=%h ctrl=%b%b%b%b%b%b out=%h zr=%b ng=%b", $time, x, y, zx, nx, zy, ny,
               f, no, out, zr, ng);
      assert (out == test_cases[i].out && zr == test_cases[i].zr && ng == test_cases[i].ng)
      else
        $error(
            "Test %0d: out=%h/%h zr=%b/%b ng=%b/%b",
            i,
            out,
            test_cases[i].out,
            zr,
            test_cases[i].zr,
            ng,
            test_cases[i].ng
        );
    end
    $display("All tests passed");
    $finish;
  end

endmodule
